// this is first ntt implementation without mondgomoery
`define NTT_OMEGA 17
module ntt (
    input  [ 2:0] in [0:255],
    output [16:0] out[0:255]
);

reg signed [11:0] dwindle [0:127] = '{
   -1044,  -758,  -359, -1517,  1493,  1422,   287,   202,
   -171,   622,  1577,   182,   962, -1202, -1474,  1468,
    573, -1325,   264,   383,  -829,  1458, -1602,  -130,
   -681,  1017,   732,   608, -1542,   411,  -205, -1571,
   1223,   652,  -552,  1015, -1293,  1491,  -282, -1544,
    516,    -8,  -320,  -666, -1618, -1162,   126,  1469,
   -853,   -90,  -271,   830,   107, -1421,  -247,  -951,
   -398,   961, -1508,  -725,   448, -1065,   677, -1275,
  -1103,   430,   555,   843, -1251,   871,  1550,   105,
    422,   587,   177,  -235,  -291,  -460,  1574,  1653,
   -246,   778,  1159,  -147,  -777,  1483,  -602,  1119,
  -1590,   644,  -872,   349,   418,   329,  -156,   -75,
    817,  1097,   603,   610,  1322, -1285, -1465,   384,
  -1215,  -136,  1218, -1335,  -874,   220, -1187, -1659,
  -1185, -1530, -1278,   794, -1510,  -854,  -870,   478,
   -108,  -308,   996,   991,   958, -1460,  1522,  1628
};


endmodule


module cooley_tookey(
  input [15:0] a,
  input [15:0] b,
  input signed [12:0] zeta,
  output [15:0] out
);

  localparam MOD = 12'd3329;
  wire [15:0] t;
  assign t = zeta * b % MOD;
endmodule
/*
0000 0001
1000 0000
*/
