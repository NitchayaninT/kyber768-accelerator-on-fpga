../src/params.vh