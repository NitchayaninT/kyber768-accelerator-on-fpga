`timescale 1ns / 1ps
`include "params.vh"

module add_tb;
  wire [`KYBER_POLY_WIDTH - 1:0] a[`KYBER_N];
  wire [`KYBER_POLY_WIDTH - 1:0] b[`KYBER_N];
  reg  [  `KYBER_POLY_WIDTH : 0] r[`KYBER_N];

  add add_uut (
      .a(a),
      .b(b),
      .r(r)
  );
  reg [(`KYBER_POLY_WIDTH * `KYBER_N) - 1:0] a_flat;
  reg [(`KYBER_POLY_WIDTH * `KYBER_N) - 1:0] b_flat;
  genvar j;
  generate
    for (j = 0; j < 256; j++) begin : g_mapping
      assign a[j] = a_flat[`KYBER_POLY_WIDTH*j+:`KYBER_POLY_WIDTH];
      assign b[j] = b_flat[`KYBER_POLY_WIDTH*j+:`KYBER_POLY_WIDTH];
    end
  endgenerate

  int i;
  initial begin
    #10;
    a_flat <= 4096'h77d87e40446092ee1d9b820409aedf30bc41377d90d495476f23e41fbc047ac8e07fe53ec100b2e9411e096c627cbf9b1640062468fcd55c018127d630fffdb1a9c57ff566da5f9284a233486acbf40a46ff1eaf4e39bcdb875d50588028396b723dbebee4ac5ef0a1d94d482057a26ac87531aef72362ff27978b76df891db50909911dc003942c581752434551147ff8b700893958f4de850b73523ddf369cc2a76b00fd532376e5ab9caaa1e146daaf473464993ef2fa0e196f86e66f45e5b7e2da57d6900a431892ffdce5f967773c475b4325855517718d7db30110c52d61bd67abed9a76611ec7b3a843099d1919bcfec76955fbd833fe7384edb323e5eb93277020d79575675f0e8eb4db41b85b837f4fd556089a1712a22aedf6c2ba52c98b9612e89bd68193620e27ef8ae8569ecc7062389cad4c8294bdc3a2d9d471811925788785f9db4d17f49f5eb3594c06bc638e4e7748a6e93449084881b0efb087d4b5844c6452ecba9a4fd9ac940bb60c83ad353325234435c341f7a2b079f956d955b41a76b72bd5c1e2ba0c3fcf4728df087d6a3130f50782a996bcbc642ea2cc46aafc0f5552e5839a76261cbcac425fd6bf7ea360ea94bd597207202f0653f0be3568e9da88ebdec1906aba2f73e0de8f51f56c7fe92fbaca6408ddd610dd4852faa8c7ce6dcba51f4d8684cf39c17eba4c6fc6158224cd754a01a3;
    b_flat <= 4096'h347a82854a2947169558c132664d47ab8994c53e4851e7db2a8efd40cd96ea8a2cefa1c4f22a95be0d1deecfa13df9c3d89c5b76a0a45905b17ddfcf0e74f98cdc129a170166eadd684e65aeb0b12a04d62b0e83668504e5a49d1ca3bfbfd0c325340c1c501a6b258bb72f76638c5df073838e6ccb04327bc6a2b80051269fe1899db9a6240f1c10390d6b113e04b69763f539c051c337d41c0468b2e29144b6d38743475852f61e13f266aff7b31f4e41acdca3597340d50e913da12df3a44a0396807b0048058b835af812c5adcc48b0ef18a86ee2a997170922d484bdeecbf7359f64714cad8effb307a87da5cc194c2bdc0cda96350245d29a5e15dabebcbf2ba5c574afa1088b18cdc1301be565521f73a7ed28961515302bb647118d740cc7187584ec6126b5df19b45c85bf4f559a92b07207504599f20249651c986a48d3d7baee4ceb204ae469d93bd7e11962380d5cfacc53cdee6eda76024b74867a9bd6bbd008c3774bd9480e7ad02bbb7871f96ca3f0bf145d2aca939f335b6544961411c4160870da450804a1b97091444707f7c9661dbddebbd88cd4b2d81057e17d8223d5c0802074c384b9902ef397cc2f6600b18fa31d8d573a2d16005b34f6903c3fdcb115bd10706cf8104173e45623a40fac324289aec50117c4592b8f9c93410c63acc37df115ee233ade78f995e449a7ab94e2bd20ad194da4f5ad;
    #10;
    a_flat <= 4096'hb8745f9929d2420576f85831bbea9177d9b31276332ad1a2e442a3677d304f3624917b6cb682fd7d619156d8c1cca3edf6309059b906eb8fdc0251996085c8f54dc5715e75e957d561239fce091a549589127866f21ab48e9299dcbe385a67bb2f98db067098195403c97bd45b663c3823d252ac9b9776ea9dc48e9a8402b60533db16c21aa6417fab60bfa2bb9ef250ae53e1067bb01e51fd11bce740d2bd83f162d14cb40b1772a6866459e9ffc27681c2998e4809625768c343aeaa8cca0403a0bea9d61ab45f44f127857bc4f8690a6c766201fe18f29173bb31bacfc135c7b85b5f12a04dff280ad56ed77b568d13ebdf502e9f741d5c874957ec98e93dd3c1220767cdceef667c8ee8d6860edd960084a37bdf29439aa9edc23d4e934bafaba87c73e8f370d34e6191a0c1d9dec5ee18768180570a7c7f152146a4521e3889f1537cfaf3d917144c08a350a5356c75860f8bf787a770e436e7d8cb7522fd468c5049f44e261de7fb1ec57381ab616a121565bdfe1d68e95dbcab89af73837d8b69c99852e0de8a5be0426797561727550c8aa2f0e1a1b3e751437394dd4f85c035863cff17453c252011c6d767f9348cbab71edac4e6895f886966d078f2b87638a077b7c0a8295d34e0cab28a870b1daa07f21f3cae99f1075a2ddc2e000b84ced5d8e85f95dba26eac1763de2a2c78cda8e9846442751152b59cc732;
    b_flat <= 4096'h6d050d5052aca832d907cd1abebb61e53b4b597599d251e4bf1b22610695c8adad4abe75012eadf609f5737561c4960302c9383d3a571272fee26a2ee1eb2cff04c3d3dd51d3eab8b9d145d14e5c778e9d7959bbfcff78f6885e723f9bb2ef8040ef923142afb74c47179445fc52e22734dffa1492eb4b7cb1fe7c839c8290b849e260a83dae8b9ae1e178d823f1b60a54f0ca19494f837886547153432b635428412e402b1191cdca5130cd4021b3a155618e06fdcfef47821905aa77d5a9a31a48d744ed414224a11f2fbba83602b9b949bb3a5ccddf8bb4086c5ab7ddef68dde06d25c8ee8d7b556025b750ef144ebab78096a87a7f198573cc575f1d8e7ebd9e381d6ed3a5aae21137d160870277591d2f44d2f4a7205fbc625159ca12b675a30f5f2859b23ce7f9e5661452aadfd5141c9dd2472678ead031ccdf2965cc83a8b359ceaa0ec88d29d7b9edaad0b26965bfc2da724607b78fb49f98c57af24d8cfa9a44958e7568f6be9d5603e1790a066694624e279fa5366f3a8920d1a7062e14621a53f736f4770fbe649d304ff705c4829ad434075c422a7f4695eb35c650b1bffde9a0c17b8717040b2534437acccdd64131c2691e20dc5a637384244dd2ea2324fdea838a89aad3b6b8d407cd010c15fa11f1bfe54e8f7b80c8a2f153591c392f2a8e19a2d60da1d9ed1af5686df5c09ff361970da21d8c6867ae8f;
    #20;
    $finish;
  end
endmodule
