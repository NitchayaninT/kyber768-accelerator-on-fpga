module ntt(
  input [2:0] in[256],
  output [11:0] out[256]
);

endmodule

module cooley_tukey();

endmodule
