`include "params.vh"

module add(
  input clk,
  input [`KYBER_N ]

);
endmodule
