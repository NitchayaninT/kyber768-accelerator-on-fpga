`timescale 1ns / 1ps
`define DELAY 3
// for noise, gen e1,e2,r in kyber768
// e1, r = output poly 3 times (1024 bits each)
// e2 = output poly 1 time
// for public matrix, gen A transpose (9 polys)
// run once, collect 7 polys?
module public_matrix_gen_tb;
  reg clk;
  reg enable;
  reg rst;
  reg [255:0] seed;
  reg public_matrix_done;
  //// output
  wire [3:0] public_matrix_poly_index;
  wire public_matrix_poly_valid;
  wire [15:0] A [0:8][0:255];
  reg [15:0] coeff;

  public_matrix_gen hash_top_uut (
        .clk(clk),
        .enable(enable),
        .rst(rst),
        .seed(seed),
        .public_matrix_done(public_matrix_done),
        .public_matrix_poly_index(public_matrix_poly_index),
        .public_matrix_poly_valid(public_matrix_poly_valid),
        .A(A)
  );
  // reverse bytes for printing (this time, per 4 bytes)
task print_decimal_pm(input [4095:0] S);
    integer b;
    localparam integer NUM_BYTES = 256;
    //reg [4095:0] reverse_coef;
    logic [15:0] coeff;
    begin
        // reverse bytes (for visualization)
        for (b = 0; b < NUM_BYTES; b = b + 1) begin
            coeff = S[16*b +: 16];
            // print as deci
            $write("%0d ", coeff);
        end
    end
endtask

wire [15:0] poly_out_debug[3][3][255];
genvar x,y,z;
generate
    for (x=0;x<3;x++) begin
        for(y=0;y<3;y++) begin
            for(z=0;z<256;z++)begin
                localparam int p = (x*3)+y;
                assign poly_out_debug[x][y][z] = hash_top_uut.A[p][z];
            end
        end
    end
endgenerate
initial begin
    $dumpfile("dump.vcd");
    $dumpvars(0, public_matrix_gen_tb);
    //$monitor(" phase:%d\n enable: %h\n index_i:%d\n index_j:%d\n state_reg: %h\n bit_squeezed :%d\n output len:%d\n output string:%h\n done:%d\n", hash_top_uut.shake128_public_matrix.phase, hash_top_uut.shake128_public_matrix.enable, hash_top_uut.shake128_public_matrix.index_i, hash_top_uut.shake128_public_matrix.index_j, hash_top_uut.shake128_public_matrix.state_reg, hash_top_uut.shake128_public_matrix.bits_squeezed, hash_top_uut.shake128_public_matrix.output_len, hash_top_uut.shake128_public_matrix.output_string, hash_top_uut.shake_pm_done);
    //$monitor("index: %d\n rej enable: %d\n, pm poly out:%h\n rej done:%h\n running:%d\n",hash_top_uut.public_matrix_poly_index,hash_top_uut.reject_sampling_module.enable, hash_top_uut.reject_sampling_module.public_matrix_poly,hash_top_uut.rej_done, hash_top_uut.reject_sampling_module.running);
    clk = 0;
    forever #(`DELAY / 2) clk = ~clk;
  end
integer i,j,k;
// for printing public matrix
integer round = 0;

reg [2:0] prev_state_reg;
/*always @(*) begin
    if (hash_top_uut.shake128_public_matrix.phase==4) begin
        $display("\n\nOutput of round %d", round);
        for(i = 0; i< 25;i++) begin
            $display("%d: %d", i, hash_top_uut.shake128_public_matrix.state_reg[i*64+:64]);
        end
        round++;
    end
end
*/
initial begin
    // -- INPUT -- //
    rst = 1;
    seed = 256'hf8f11229044dfea54ddc214aaa439e7ea06b9b4ede8a3e3f6dfef500c9665598;
    enable = 0;

    // Release reset to start loading state_reg, done, etc
    #(`DELAY) rst = 0;
    #(`DELAY) enable = 1;

    //wait (noise_done == 1'b1);
    wait (public_matrix_done == 1'b1);

    #(`DELAY * 10);

    for (j = 0; j < 9; j++) begin
        $display("=== Poly %0d ===", j);
        for (i = 0; i < 256; i++) begin
            // pack 16 unpacked bits into a packed vector
            coeff = A[j][i];
            $write("%0d ", coeff);
            if ((i % 16) == 15) $write("\n");
        end
        $write("\n");
    end

 end
endmodule

// CHECKING PUBLIC MATRIX OUTPUT
// Public Matrix from SHAKE : b17a22ce5d458ba33d6931d893324e04123b1590846653d49d019a59da9ddd1aad293fc43863b0f63c093b2e9325249a0e45cf390f8ea91fdf9450a90c34babde106958e80184c9dfcf78da5f66fd7f65feef73aced58d4d995606c2ab56d11141ec5e47c6c8baaa5fcc346f9ea76c58389af2cf4df93f38c70f542cbae644577d22fd10d46f4f5c70d72c99775bc9ed7e0c417b6af0e9e545603f42df15d09481539cfef0bdb84b3899339793c2759f4c6d3b73f07f5a2ef7927f39a6ca2b45102a5b2794449c99b04617b2bee4777e043007a9e07eb858f4a49fdb5380e1de3b739c795715f4fc11223f37896d5fce01f63ce25780c462a6f9379a8d112d026133e5b6b6df3795cc374c51785f435d2bcf64e4f6be21e38f7d8c1c447b2e73b9ca12d58a71efbc7d4cae4cb99541d8f5662dc2ad1b4083c449461b60e7ca6bd395bc878cd37eff6ebca7ec10ee6ffbe1f719eec9ebbfd31e60b174c4e4a2940d14ce9343b3c10d9ddd42d92d04c19c1ae1901cb4095fa4e00ee14949ad2f513257e1bc6295e8a0eda314c3ac3b67a0d62a4397efedd96eed0ecba9cc195276800fa0bd99a52dcdbe8d959276e5ace0fb215f3a7b01d781ef77287786653a6e7a15c187709b16854e142910976b0987ac13fd54981c47af0635eb286caeadd9c25c425088160c7965659c1e659c9a5942b330dd5f045ddf6689eac9ea06a1bd59b27768331e8b8d74f8b5c661789989160286a71e740bcd0718d5e8b84a05bdb9aa0964512c452e2feec81ad94069ce5430a05d5b806d311a9a913492a419012859b1884f94698c62a85ac0d7cf91e370d3a14a0d75d1ee3177b29cdf4aac5463b73d722603fcd1c946b71f4d60b1d0619be63b2c10464e8eed2db46d0fa6ba16beaa63a2f5f9ff6ccbe3e70953c633e81da07d3389ef6becfcfdba740b56bc
// After Sampling Rejection : 07100291044e0851069b070807c101570a6e03a605860772087701d700170b3a05f201fb0ce50769029508db02da05990bda000f08070652019c0ca90cb006ed09ed074302ad06a006730bac0c3104a300e8095602bc07320512049409e100ee00a405f009b401c900e101a90cc10042042d00dc01b3043903ce01400a2e04c4074b016001ed03bf09ee019f07e1010e0ca70bc607ed038c087b0c950bca001b046409c40834001b0adc022d066f05d8041905b904ca07db0cef07180ad5012c0ab9073204410c8c07d8021b04cf02b505f7085104c307cc095307df0b6b06e50336010202d1018d09a307f90a6602c4080507e203cf06010ce50893073f022101fc055707990c7303bd080503db09fa04f4058b087e09070300047e077e04be0b2107460b09099c0449042705b20a1004520bca0a63097f092f072e05a707330b6d04c90c2903970339093804bb08bd0538019405df0423045e05e90a7b04100c7e095b0779092c005c04f6010f07d507440a2c0540038304dc09a3085806ca079e06f304cc05fa0aba0c8c064705ee0c41011d01560abc02060569094d08dd05ce03af07ee05ff06d706ff06a508df07fc09d40c180808006e01bd0ba3040c0a95009408e00cf4050e09a20425093200930cf60b0603380c430ad10add09dd0a5909a0019d03660849001503b1020404e30293016903da038b045502270ab1
// Reverse coeffs to compare with C : 0ab102270455038b03da0169029304e3020403b1001508490366019d09a00a5909dd0add0ad10c4303380b060cf600930932042509a2050e0cf408e000940a95040c0ba301bd006e08080c1809d407fc08df06a506ff06d705ff07ee03af05ce08dd094d056902060abc0156011d0c4105ee06470c8c0aba05fa04cc06f3079e06ca085809a304dc038305400a2c074407d5010f04f6005c092c0779095b0c7e04100a7b05e9045e042305df0194053808bd04bb0938033903970c2904c90b6d073305a7072e092f097f0a630bca04520a1005b204270449099c0b0907460b2104be077e047e03000907087e058b04f409fa03db080503bd0c730799055701fc0221073f08930ce5060103cf07e2080502c40a6607f909a3018d02d10102033606e50b6b07df095307cc04c3085105f702b504cf021b07d80c8c044107320ab9012c0ad507180cef07db04ca05b9041905d8066f022d0adc001b083409c40464001b0bca0c95087b038c07ed0bc60ca7010e07e1019f09ee03bf01ed0160074b04c40a2e014003ce043901b300dc042d00420cc101a900e101c909b405f000a400ee09e104940512073202bc095600e804a30c310bac067306a002ad074309ed06ed0cb00ca9019c06520807000f0bda059902da08db029507690ce501fb05f20b3a001701d708770772058603a60a6e015707c10708069b0851044e02910710
// Coef from LSB to MSB order : 2737 551 1109 907 986 361 659 1251 516 945 21 2121 870 413 2464 2649 2525 2781 2769 3139 824 2822 3318 147 2354 1061 2466 1294 3316 2272 148 2709 1036 2979 445 110 2056 3096 2516 2044 2271 1701 1791 1751 1535 2030 943 1486 2269 2381 1385 518 2748 342 285 3137 1518 1607 3212 2746 1530 1228 1779 1950 1738 2136 2467 1244 899 1344 2604 1860 2005 271 1270 92 2348 1913 2395 3198 1040 2683 1513 1118 1059 1503 404 1336 2237 1211 2360 825 919 3113 1225 2925 1843 1447 1838 2351 2431 2659 3018 1106 2576 1458 1063 1097 2460 2825 1862 2849 1214 1918 1150 768 2311 2174 1419 1268 2554 987 2053 957 3187 1945 1367 508 545 1855 2195 3301 1537 975 2018 2053 708 2662 2041 2467 397 721 258 822 1765 2923 2015 2387 1996 1219 2129 1527 693 1231 539 2008 3212 1089 1842 2745 300 2773 1816 3311 2011 1226 1465 1049 1496 1647 557 2780 27 2100 2500 1124 27 3018 3221 2171 908 2029 3014 3239 270 2017 415 2542 959 493 352 1867 1220 2606 320 974 1081 435 220 1069 66 3265 425 225 457 2484 1520 164 238 2529 1172 1298 1842 700 2390 232 1187 3121 2988 1651 1696 685 1859 2541 1773 3248 3241 412 1618 2055 15 3034 1433 730 2267 661 1897 3301 507 1522 2874 23 471 2167 1906 1414 934 2670 343 1985 1800 1691 2129 1102 657 1808
// From C official : 2737 551 1109 907 986 361 659 1251 516 945 21 2121 870 413 2464 2649 2525 2781 2769 3139 824 2822 3318 147 2354 1061 2466 1294 3316 2272 148 2709 1036 2979 445 110 2056 3096 2516 2044 2271 1701 1791 1751 1535 2030 943 1486 2269 2381 1385 518 2748 342 285 3137 1518 1607 3212 2746 1530 1228 1779 1950 1738 2136 2467 1244 899 1344 2604 1860 2005 271 1270 92 2348 1913 2395 3198 1040 2683 1513 1118 1059 1503 404 1336 2237 1211 2360 825 919 3113 1225 2925 1843 1447 1838 2351 2431 2659 3018 1106 2576 1458 1063 1097 2460 2825 1862 2849 1214 1918 1150 768 2311 2174 1419 1268 2554 987 2053 957 3187 1945 1367 508 545 1855 2195 3301 1537 975 2018 2053 708 2662 2041 2467 397 721 258 822 1765 2923 2015 2387 1996 1219 2129 1527 693 1231 539 2008 3212 1089 1842 2745 300 2773 1816 3311 2011 1226 1465 1049 1496 1647 557 2780 27 2100 2500 1124 27 3018 3221 2171 908 2029 3014 3239 270 2017 415 2542 959 493 352 1867 1220 2606 320 974 1081 435 220 1069 66 3265 425 225 457 2484 1520 164 238 2529 1172 1298 1842 700 2390 232 1187 3121 2988 1651 1696 685 1859 2541 1773 3248 3241 412 1618 2055 15 3034 1433 730 2267 661 1897 3301 507 1522 2874 23 471 2167 1906 1414 934 2670 343 1985 1800 1691 2129 1102 657 1808
// Reverse Sampling Verfied : 16/1/26

// CHECKING NOISE OUTPUT
// Noise from SHAKE : 99abf40515a7387aa7a41f83840467aaba58818583cae85ec7710efbeb5dce0a5e91f3fa854b8570aaa4393e663ef90458d0d9823e682c1062947b54c496ef8a9bb38198777295bb264c790628226b8a3a3ce2172d0d0c5534d8dc67d0c1155c4a98b3559c84fa82d90e4cfc474b2fda6b38ca4f0ef964bd4efd4b5cd5be6696
// After cbd :  00000000000000000001ffffffff00000000fffeffff00010000ffffffffffff0001ffff0000ffff000000000000ffffffff0000fffe00000002ffff00000001ffff000000010000ffff0001ffff00010000fffefffffffe0000ffffffff0000ffff000100000000ffffffff0000fffe00000000000100020000ffffffff00000000fffe00010000fffe0001ffff000000000001fffffffeffffffff0002ffff000000000000fffe0000ffff0001ffff00010001ffff00010002fffe00020000ffff000000000001000100010001ffff0000000000010000fffffffe00010000000100010000000000010001000100010000ffffffff00010001000200000001ffff0000ffff000000000000fffeffff0000ffff000100010000ffff00000001000100000001fffe0000ffff0002ffffffff0001ffff0000ffff00000000ffff0000ffff000000000002ffff000000000002ffff000200000000ffff0000000000010000ffff0000ffff0001ffff00000000000000000002000000010000ffff00000000fffeffff0000ffffffff0001000000010000ffff00010001fffe00010000fffffffffffffffe0000ffff0002ffff0000ffff00010000ffff0001000000000000000000010000ffffffffffffffff0002000100000000ffff00000001000100000002ffff0000000100010000000000000000ffff0000000100000000
// Coef from LSB to MSB order : 0 0 1 0 -1 0 0 0 0 1 1 0 -1 2 0 1 1 0 -1 0 0 1 2 -1 -1 -1 -1 0 1 0 0 0 0 1 -1 0 1 -1 0 -1 2 -1 0 -2 -1 -1 -1 0 1 -2 1 1 -1 0 1 0 1 -1 -1 0 -1 -2 0 0 -1 0 1 0 2 0 0 0 0 -1 1 -1 0 -1 0 1 0 0 -1 0 0 2 -1 2 0 0 -1 2 0 0 -1 0 -1 0 0 -1 0 -1 1 -1 -1 2 -1 0 -2 1 0 1 1 0 -1 0 1 1 -1 0 -1 -2 0 0 0 -1 0 -1 1 0 2 1 1 -1 -1 0 1 1 1 1 0 0 1 1 0 1 -2 -1 0 1 0 0 -1 1 1 1 1 0 0 -1 0 2 -2 2 1 -1 1 1 -1 1 -1 0 -2 0 0 0 -1 2 -1 -1 -2 -1 1 0 0 -1 1 -2 0 1 -2 0 0 -1 -1 0 2 1 0 0 -2 0 -1 -1 0 0 1 -1 0 -1 -1 0 -2 -1 -2 0 1 -1 1 -1 0 1 0 -1 1 0 -1 2 0 -2 0 -1 -1 0 0 0 -1 0 -1 1 -1 -1 -1 0 1 -1 -2 0 0 -1 -1 1 0 0 0 0 
// From C official : 0 0 1 0 -1 0 0 0 0 1 1 0 -1 2 0 1 1 0 -1 0 0 1 2 -1 -1 -1 -1 0 1 0 0 0 0 1 -1 0 1 -1 0 -1 2 -1 0 -2 -1 -1 -1 0 1 -2 1 1 -1 0 1 0 1 -1 -1 0 -1 -2 0 0 -1 0 1 0 2 0 0 0 0 -1 1 -1 0 -1 0 1 0 0 -1 0 0 2 -1 2 0 0 -1 2 0 0 -1 0 -1 0 0 -1 0 -1 1 -1 -1 2 -1 0 -2 1 0 1 1 0 -1 0 1 1 -1 0 -1 -2 0 0 0 -1 0 -1 1 0 2 1 1 -1 -1 0 1 1 1 1 0 0 1 1 0 1 -2 -1 0 1 0 0 -1 1 1 1 1 0 0 -1 0 2 -2 2 1 -1 1 1 -1 1 -1 0 -2 0 0 0 -1 2 -1 -1 -2 -1 1 0 0 -1 1 -2 0 1 -2 0 0 -1 -1 0 2 1 0 0 -2 0 -1 -1 0 0 1 -1 0 -1 -1 0 -2 -1 -2 0 1 -1 1 -1 0 1 0 -1 1 0 -1 2 0 -2 0 -1 -1 0 0 0 -1 0 -1 1 -1 -1 -1 0 1 -1 -2 0 0 -1 -1 1 0 0 0 0
// CBD verified : 16/1/26

// Public Matrix Streams from SHAKE
/*
1.dbe65936fac169bd5d7888e1012ca9df90cb3392ca34000e5fbaad4c95d06f27664952e488193d313722ca38591337989f502d9188faafb9b9472b6d5c85948abb752c72483f54a2bd80378740052ddcd10e55b9499f0ec1ae2487b6931fbefd29953a7eaa0d36a614812dbb8466036a0866b98c2740b864c8a679f051599c8667b230bd85ccbd294e7f3d7c2edfc9532d47791f77e0aff4425da8199b48eb9e3a44b40d24ce21f19d9747aa41c3ca9a0f40b4a8c79e1bdaf86fb52cc226373fa523bab2af1e46e5fd046f4dfd05137d5dde7c1bcb584e717e93d03e8f9d1a4a8bf581f7455d44f4dc0d8e25913e82c417ef29bf2d26cddac2c9adb74efeeee4e6d3f13faaa12e430258e5c7a37c37584db6fab6008f8832003b15d0a5af18dcc766496b922242012a8a2a4c0511ac71476629fc9d5871939278803bdf9ec049e75f83da4956fc4e7c9b62307e6ffdf1a73387ae69ca267e8cd9844473bfc24ce6b08ab9447dca14a62a032514b71a3d69f3e532152c68d02180c170ca99951a748a17592011d946dbe3e0d14d8e4005e90c19189ff2826a94a067ac021ac76db1699ee2b6ddda083f45e29e2d537e4500032536668d5917fb1c4fe8a73f31799a3df8b130d368513b3a18a24f6623207337249b137851d67624c458ce6cef1a63257e3d92cb61cce10f9e979049a6d9b3194fcaa2f5743b976a9de7b4dcf61568e639cf61df867ba391d6f27bca44f5adac07e09e088cda63f8a5214450ce313e350c10a65d34975041a73f78c8968c6e75a0895adc506359095ccdb936cbbf2426fb53fdc53414cddeb8d6a95de8a9debd8634ebeb861ca0d3551feef5f4b39154acb90c697ec1d25101950fac0623a53fef8647ce485b07a082e9c2d7dd598b053984b21916ee66a153528fb631255541f9b4e5ae8fe837a706c2ced50679
2.f267fe4749667765c0109c2004dc7b070c695b0fabbcfb0d190f71fbd1e2420f4bfd97ce6d2868b3445840f0ec93f058639dcac9601e0786eae28b69b884b650e9caa1ea417c13388235ac4c68c20f24b7b3da6e00ddaeb5aba79861f0f46bc57faaced94bc8e49d958bab9165f2c2850edcee5861583c02d01c8a712a86df231a718da7702403678fb61adee6565cd58b4fac0a7e9ecc4c541ea89530091015c85f73a14ffa9f8ff30e4bad549d34d51d133682ef8dec0964f01e15127ef38c12510ff5ad546cd6480cd7eedfa73177301edf1e434cf2deaab84bb63eb98a971e0e595cbc4ce956e18e6613b6da2057f3a0c103c7bab1ec19ea212928554baafd2889fb6b3c0d0b816d7f2732d0754a953e5f14d5c1deb4b3fbdb93368a1469b9c62aba3d82809a90138656346bd1d672bb742f648d2a5a9c9a8de873c3bbabd737136c8a8aa97e6b4800883c470e039fdc2670754b7ce6d446b8a017f161ce6051af635dcabfa14a487c7a57f86843cafaa7ff420c6a63c80ad9bbc4d58d15eee8dbf3e3b21de103a64fa142909e4d4b620de55790df390b4e3eaaf0efa2d4e0b1a5e671b2cae6fb50002d5e88e1646197d43df25759aa1f17a19c08c1172ba5e7b9e8aac89b2172feeeda13c62fa0e0d46c2776439fdcb6a0f75ac1503b60ee08100cd350ca5a0e3361d3da832ac2ec9df323c31bb59084dc8d21a492af8497ffc1cf4d1ea016ce787b09c9c4825adf29cc58e0ee124d7e5d24f444868af39c63d647820679f1ae1a93ea7b3a305e1f2bb6ebc72034b472511c1e75c0447f83f75b1cbbd7795c7f6b81bc6b369588e812cf0ed06de21a876755dbaa2d097fa473ed08eb850107fe3ed04c7e92bad14df79900bd36352b007f66ce887697d3aab8f7b0487c6523808b12348640318d0250d0caa7cfb320bafe28bf7a3442ed
3.a798ead47cd0d0de2fb67565627517a36640432d45eaa698abd1a9d9fa34800d56fb5e33eda694c5b9884f575eeea3c076f0162e9adf3c4f4bc000103a81f69b43c68e8b0be2df84442fc9e8ae2369462f233f51953f3b6dbb50abce148626fd2bafe2d33572becd149610c931c426dbe29408e5560c657a59faa002f4a39f651f5317169a6209e9f2d03f6c1f26f72b5adfaa2f1df3f551ddbf4f6030c3cf69fe3fc3011ff3019fbe84124f9498b778728fad0066c71b3f8b0ec1d8e19f5ac63f9ef6ed943b12d4a7e3ae7beaea04a4deaab48ac8f977c9ce77fc4676024507056765d1a3bb03f4063e5f1a5b11bc55ee166c58338bc2f3dde96ac5d77fbe5a09f31e08b880fa495c21ca5280fd09e52652e771c098d073014630237df35eb18aa8a5593bd1cbebf120064847f4ffe630945cfcbe0d6ebec9b8273a56b516883c6ba36d0437e344167eb023ec32e1b1fa257fef0e3fe4c07bcf2030119525ec63e0151e36f1950cab4d2c7504f631ed5f62adc120c0f330d536deaa1a796f9eaadb720729f9a9f06aeb4875bbe740f52e636c54d9ed35cd17085dc010f7f34ec3eae43c37bb09583c4b6f67879cf95cac0a81281eeffe07f1270bb7601afb0077df8231f2857901269dc345b583326fd1dab7c1d1c1b00cb5cd2a62ab72674308744983f85dd4e4ddef4ecb9299dd9bf932b3262998bd4797ac765363cdde040f18e759331ad9e26713cf153761075429413c87e0d55f0170bb41a57c9e66a94dbdb04bc523db9f46e02871f4d9b6955b7d015bd66144c30a4c50da63dc0b8d8b1572302f9b17ea3f212cc6f2354ff854c35a0520abdb6bab70b35de5edff5adc61c4d8af7bff34ab562734054b2926b256de63f5591d97f94cb3b75222eaa257f2f0c1aa4180d2a3bdfd96903eb6ae8324ff18982ba19abef0908131472c12
4.6755eca382f34f3e9b7b26f67de864f5fae38f9c0d154fe958fea5d75e50feb920f8f47a18a657ecb14da08a5e20b9233dccbca657f10b8ac18da670a9e1bd0b7c4b7ab68e217d203084f51e81a46c4dff96a99c059ca502b177b8f0b9e2dc9b944b1772e980a1057b216c3d5696a2bf05fcbaf3e04e757cc7aa0ac156f20535848092de5f5dcf1e38c0ca1a7f4795da8c7e9afd4c1d8cab3243edd99c527b82b6d41942788b1d2e39908023d4d7ec1a1b189c54ada8fdcef8b2b6f1bb68a41e3121328cde57f0fd175a4c508356a4b538c3df1de1b631746a14baaf21bb3640e85bd6763dc12ccee40120f8ff769cea481d0775dd0f3950c5794fe745b85b6e4bec543a7314ad89281754124349cb13a1bc163d7514ecf76700206faaef610deecefb71c5cf02e0c8bbb4dd23207b48b87266cc890a84c0e0d3f21cb0418de24e926539f1a5ab270032fec7047764d454088134ae51be6e2a639caca9e6a09d4349dc781a4316b399513ef078e8a20a8610342cfbe1871401c0acbc9c5468c90dc84e3ddf1f99896a7437188492a512427b344d97e555df97c4b8af69a2ce059654cbb4ab78e6c54784cbef0046b615a124de2e9f2eef40686a299f54e2adbbfb97548fd3fcae5e07fcd84ebab4ebabf1838a967bb0e7f495528e96c9a4d18ceda3b95a48943fab108dac099218c96484405c77300b40ad9bbdaa0361b7fc292ba06e7c16215aac89eff58d91430d86d55e67cc7722a523ba25cfd1c37d11b70480517062cb1c0b6738dcb81ce120a56e8e3d75849fd6b70d55b57fe9c98c22956a21aaaf048d4fa54a3de517cd4eef46023b427b586bb7e7b50460dd215591ed861f50a090ae3da9d998843204a585ddf8fd9c059bf0edd2225b5d39649019b45ce8d34af6a9e7f24ae44cc27a68b5482826d81258991dfb4113b030af8489
5.93569dcc08da6997c8f376c8a65b479c710d06aec45177544a950ecfa59d4a26aec77598d27f56a555532e41e5e034c8ec13327706c737f5a49b9249d31c699c3daf539a995d5d8ed548074b40e366959cec6df843fb3682cbee16c4af99c0098dcdf1dfb8b1c4f980d42a554c44c084ba3b405fa3edda75d8f07a26f6e999b4b0170203c579deb3ce677df5b302c4e6cf8b10355163fb9e25102d452a72ff481c97574c058438d15470db7d371afab6bdc1ca629581a99d315beb6f7ad2f12045082316a9fb4f7fc6077ed21d126fa857582152a57564f1a019a93be7f03c25fab66a5777d3031e1365e7116c84291c2882a3c97eb85b2fc04492779ae8128fa2a88c45675fa77aaac8af4390c3891b611b453b5533e89c3fdf917fe440cf829728e6bf783e6354a220387b7c444915621f9d997978d2e74861fff3562932d326b306eacba88e9cc15ee58f907721ece58e8ef8b7d49083d01f6db23e1be888ed194821833da353b9a163a2ed8b444d685157fc35a9661628929d207fbe7dce4f4720e88014a00c635355ab26fe56d9b41d9b461edc16042391b1e57eba08c462f6eb19a650987f366ae905eee68116bfdadcf90b584ac582ac4d5307aee60e5cb65cda6d1fd4c78867fe8d666953bc309fdef4ac97692bb2625a0b45ed0aea744444b7fbdb86a76767dfef99889ae39fde1a5209d501418fe741c6d5679f419e5010679f26c8bcd193b15e15de452528c25df45077df7dfea03e13c153ceed74e9c4256ff8056def92676dfb07c5951a823020f2a88645a72924e38e759e6c1725ac72da2dc3a5a7c7bacdd1f215efc92494804d0691a3e240e9d2ffa3f80798a0f6c1b723ce7b52c8176d36b3b2379c23ed17bd909524837db48535becbc881d51514d4fbdaf97e62a455c8d2dfa577ae76b16fcd40a14a415a5b73d3ce92
6.6b5af57f100149491cf321eeef197cc3bdc6728a499f7e1eb6dc4e1a920cf545a5ed9a63d1b42ef0284565373b744e3559e4e0acd508ddf9fe6bbcae05e3233882fd118fae965b6fe24cb40edc17644692f0e671a0e772ef5abbc6edf8a3ab46d0594fc09a6a56747cb64f7579cfa2b9ec8010a39b9a0bde043d3b1adda914b26c74ad3664f29d0c329993dd13b20d200eb5d70aa3bc2fc852f9500978cc4348a055d71629ab1d1dcfb78d4c088a0e1aa4b5f4a0706ae4186539be16cff43be8f69994cae1f65f4e51bf607b38fb56ca3156212cf64693809b0405d6e6927d4416623be6b8ef4d8d1e60581945e64ae4a97ae320e2d76d5dfcd64a717f0ecd677720bb62cc874ccb62df00aa15b13023aad68f3286c0c9765ff3b3c58c1f0bcd63126923deb92d26c67bcb35a2d311a1c5246e1b0885e687501e2c054f157d2afaa59c824db2771bf2b07aca1b5e003e4941d1cf7eb7a7eea3059b6c7326b9286aa8b8c6197299a717c72c5116df65089732cfb45ad7a5b4286671e8e935ffcfb5563f40fd4801d0436c014ad0f03112735c1d77dd0c1cc73d90c75c2e5c991c747292d1e214de0358a95a31edefe15b3d4ea5685e6526e97cf81431e0999ded2b2f8bcf74645d3fe8928744258ab3afacd9bc1e85ef761406e094683b132616fc516821b9c8a2c8b10fb53b354721392cf931180ea6b0d96cd81bbb8616d1c1a2916943ec1c173659f260614cab4aec5e037984dba450bc7724f19a67c4bc45376efd6ec7d1e260cad19fa312251655ff57a08cfc1f369811c1bcfefc481829804761a4cd18b0eca1de7257c5020fd57499478cd7e0a4271b78a62e3c86f6f6454a79ac01a86b707e11055695ee549325ef1ce6742030e5df02504f215972a66cce3c1e42b43065bfa26a1f2c18e4ccfca47ca6f58e584a577c26e5567f2102
7.ea13b543f67f2a90daa3c4469cc644951a9893d0a605914739de43762a853501478b2200ff3014e9cbf6c651b91a7430d4b1c7e9e52798f3b358c5f6ad8540ad0f15c88542e5121ebc779843ecd94218ed19181cb9f2bb40e3f14c5b7b07cf47b8f7c538e1cd091644cd1456e4ce2429e75ce4c25fd8aad27ffbfd84081f2864473f9e1e1d83e1d47794fcf2b98c81296e9f5d085366f873cf80512a50847b33c0bfb69814beeff65f885933910a698fbedcabf191b11656a4d7cd7b74bb0242e853f5f9b69060a9b585f35e11380da2e388decf59cf7f4f5479fcb77e1f7829973d661c1e958f3fca2e1e16b0636f0e3fab8ef22f3c8bfe90752047415f94d5c4368e1c6ef14a7597187c77825c1d56cc9fb8de1ea2a71a3f30d2697d2789c8e9fbdd897d14dd1a18f49e1c8554fda42a5f5ae5a0a949d9ba707bbf97292aa21a1492c312f8bd43148ca287e8af76610b9ff852ef165db92b4dac471c8c7db4f15c563ac59d713be94c8af878ad2d9a4b141d06bb06bf4b8403cb84450fd32854da847301e969c7ff7ca60711d7a621adddbd1eb1aec816c8a22f9809e99cc97b29481866f13efa191d9cc3f733109b860f1eea236479618401bcb47efbbf0fe8563f124e7574ff56def4efa14efaf5b15dfe4cc6d4f8455dd17862f965bdec944aa54c0c06089ba029d0c64f3f2456b7c7b1db21c8a01366a995be05ff7c4a4e6597e56995089fc70e6707e51299af575fa91f74225ee8990a013419faea61c13b11babb7285736d79ba4e70da47a7fdef58a75e0a540f39557bd95c96cd63112ff5ce90aba9ebb22580398c23dc4eb895d5d1502893a3bb98655e2ee3e6c0e63b067d74dc3ade32222c2ef446992494ee133747a53ffcad7e9df04ac4b594a7e90330d728ee8d405e4251ea619f769a82dea463a1c4d262218d90c4d1eeba
8.af6c46506c7eb910f775ea3f63d96aef64f49d4e6945782c47ad9d38b09d34198d69c974ca36210344c2bf7757e46aaa88f8998e1041893882750c1894436edaf484092dcc57fe0f08d43b461a90bfc732ee3e1dfb70174f1ed25093444550b178a8900da43833056e9596a19e91c3d557295cf5310d59e63f4943f013b2b41a274ac39e4eec2e2dc4bdf2083d5464dac871a2d8ad03f3f36588a5726afd1790f7be0ce15f63693c376cfbdfd9198ac4c091f0215e34f6f67c1fa78ddb1b2ca0bc84adcdff0730723ed99ba52252488e2fabb832052e34741febf8b486a2ce9c29d84781de813a40d705ff0e2a885be7d63c328424fcfc212cc25b3105c7170dce81cd344e025bef01f87689c9f377e355987725a84df9e8f0b76c695f07b5f8ac2946a1444311c6ea9debb37d624dc6d7439a9d5278e8687f241b9f14286e3a566aaa12026a0a68e6297a47641600ce378ac44ab8ea963ad69c40326c06662ddb077299a34ee0287be1564c9bc97ac4dd2ce5708c6d781dc2cb52f601721634f71cc048b334fb70c8f209d278c0b6c04f8840e5c4c1e02791078494f1c9032654e61f01f49e689dcd315ed3859ca756c7b73f6987e700985e163a195cde3df88a1c57112e737858828d1b1e7e785825d531d0a800e1b636da480eabd25433e6aabb21a23ccecd30eb1391186a1b2d9e745d3d8e45b01bf68e67a945aa39feea18a1751d3be4e739f9a4417015145aca08d8efc994a4fbc699c5024a2a0bab76955a4e086ae6909bb7335af1e40b0af337befd8c43c6bfc464ba11f2ac08850c5f98fc4d73697003e6d9f79c68bec44c17b1277eb726ca1aaa55ce953041a8ce161bcb993f82a27cd79a74434b65e4544ca98f2b63ae0d36157d32dfe44accef9960d524f3a0d9cc3a2dbcd750a0bd42ec93dc590a4d89ecf807e80b3ea6db3a
9.7f6008ec8e50de3752d3ed3ec7a332cb5f00957b44f8a34d45ac1acf765e02e56f7954751240deb4b2e0f8f99f024e0421dcadf16a930f2209411f897bd44fc64ec420b9fc16eaa52d988eb04a3e8e57a7f169f446c2bfa1d18c10eb834135cef8462b3882a15c7c7237bc746380e81b9e48df277f381d19f9526d62ff59e713dd460e43f799f76d9006b640e39d2f9045a69e2fd770b89052245fdfc6af5fb7d85694b5d94a34ea69b564620ccd0ea765667bafa259bebaaf78335281ccba06b0b10577737f3235d45f040541c3d99258f1427845be273b584ba1a204d7263e76c496496f109ab274a2ff98ae130da85530d3cf46b1001d93b5ccd06a13f43b5de636cba2e357e2431854f5ea4feac148adf001f06082a373122c6799443cd2c062568e67b0b9b93bad65b7a247793d9e41ae1715cf17f6873f910673e42b65669dac8e386acd1af189ed7d047b6b17e51140c17dca0a2aa024f1cb2de02ffbd41e760405624a2cdb32369154902e695e1c18a8b3750903f1a7547006be290562c86a6f4984e2185bdc715196e5cc30729a189a67b2adb1eca95023ca43a1103db4590b787644d90703772b362c26042e3e762d1a07d2f5651ca642ac8d1e0543bb818fd3cbc90a30d0082ac0e94dd45923c517ff63e47a7163af13a7cc6cba549ae83a44a81067a621542de5556c246ec570a2a45290f7bec61a75b377a6b30b9d2a652808b425609b63b9663c5c71170908e5759875630cb4405ed1ff347d4f2bd2313f5779e808e992497ed218a40516181f87f9c71f94d69523a895fe0d872a8c2f98e1940e677511420175fb8f3b095a884bb174c50cf93f1eb1a72e8af085a8d6d9b7868a41f974f7d3dc585aed96dcd9f335fd35a7aad72b0f7563a40b555c5f89992ff99a04689af7b885b4716e2d4ab6f28614edd6d96775a8e5c5
*/

// Public Matrix Poly (4096 bits)
/*
1.01ae0ce508c4024706d60517081309b2043707320023066401830a3b051608d3030b01f803d90a790313075908d6063602500300045702d904530b1601a002ac067a009406a802f209f1081900ce0905040800e306d90112005901780a7401a905990ca700c1080201d006820c15032e05f306930b71042500320aa6014c0a7d044b098a0b0e064c0c2b044804d908c70ca609ae087303a707e3006209b70c4e0649035f09c009ed080708920937015809df0c29066407710ac1010504c20a8a02a001420229026b049606c708af0a5d001503b0003208880b6f0ab604d5083707ca03c7080204320aa306e40b7a0c2d0acd0262029e0c48023e0912058e00dd0cf4044501f508b40a1a09d8037e07140cb10b7c013005fd04d6054601ea0ba203a503f307260c220cb506ff08da01b90a8b044000f90aca0c3401aa0479079d01ce024004430a9e089b019a085d042f04af071f0794072d053c09df02e70c3d07f40bdc0c850bd300b20678069c059501f0079a06c8064b084002780cb90660086a003606840bb2014a063600da0a7e03a90529093b0687024a00e90b95050e0c2d00540087037800bd0a25043f0487022c075b0b8a0948055c06d20b470b9b09af089102d5009f09830713059308ca0223073103d1098802490662076f054c0adb0a5f00e000340ca902330cb900df0a920c01087805db0c1f0a36059e06db
2.06dc09f4037602760cd4002f0c6103da02190bc80aae08b9052b017c010809ca011701fa0a59057f023d0761064e018805e20d00050f0be60cab027105b104a200aa03e4039d057e050d06240b4d09e900420a14003e011d0b2e03f308ee01580c4b0bd900ac086306a00c4207fa0ca40368077a07c4084a0a1b05d603af051600ce061f01170a0b0846067c04b70570026d0c9f003003c8080004860b7e0a980a8a06c103370bbb0c3703e808d90a9c05a20a8d06420bb702d60b340568061309090a80082302ac06b90691048a036903db03b401d5014509540a75022707f600b006bf0b89028f04b50528029201ea019e0cb10bac07030c1a00f3057200da0b61036608ee01560cbc05c5090e01e9078a0b9304bb08aa024c043101e30077031a07df070c048d066c054a00f5011208cf037e0121051e04090823061301dd053409d504ad04b008f904fa017305fc081501000930095a081e05440ccc09e70ac40c560b68003204700a7801a203df08620a7108a10cd000230c58061508ee0c2f0265091a0b8b09590c840bd90cea0a7f0c560bf401980a7a0bb50aed0d0006ed0ab30b72040f0c26084c0ac305820381037c041e0aa10cae09500b6804b806980be2060701e600c90ca9058f00930040058404b30682086d0ce907fd04b001fb071000df0bbc0ab006900c0707bd0c0402090c100c0605770664094707f2
3.04d405df088304970408043607720ab6022a0cdb050c0b0c01d10c1b07da083b05450c3900170985018207000a600b700b2707fe08100aac05cf099c0876076f04b30c58009b0b3703ce04ea0c3400c005d008170cd305ed046c0632040e07bb075408eb06af00a90907072d0baa09e601aa0ade036d053000200c1a05fe047502c400c905f1036103ec02590511030200cf07bc00e403f007f205fa0b1e013203b007e10644070406da036b03c808160b55063a027b08c90be60bef0c5c094300e60447048006200bcb0b590a5a088a0b1507d203300460017308c0071e0752026e050900520ca2015c049f0a800b80081e095a0be70c560ae903c208b3035806c106ee055b0c1105b10a5f03e006f4003b0ba30567005007450027064607ce0c9707f90c880ab40aad004e0aea07ba0a7d041203b904ed0c650a9f08c100e80b3f01bc0766000a072708b70989044f012804be09f001f301f001c303ff0cfc0330060401f50aad02bf072601f60c3f02e90096029a0161075301f6059f0a3f04020a0f0a5907a6050c056e0508094e02db026c04310c910096014c072305d30686014c050b0b6d03b3051302f40669023a0c92084d00b80b8e0c64039b013a010000c004b40a2e016f00760c0a03ee05e5074f088b09c5094a06ed03350560034f0ad90a9d01ab098a06ea0452040606a301770562065705b602fd0cd408a7
4.01a40c99068e052905f4007b09680a830beb0b4b0a4e0c0705ea097f0bbb0ade025409f2096a068400ef02e904a1015b0646000e084407c508ab0b4c0b54096005ce0a2609af0b8c049705e5097407b402120a5902840183077406a8099901fd04ec080d0c96085409cb0cac0c000114087e01fb02c3041008600aa208f003e501990b31064301a708dc0494039d0a0e06a90ac90c6302a6051a081008540477004c07fe032000270aba05f10396059204ee028d041b001c03e00c08040a089c0c66072b084807b2002304bb0c8e00020cfc057100d601ef0aa6000607f7047503d106bc0a1103cb0494031205410728089a07330a540b6e05bb08450c55003900fd00710c760820001e04ce02cc013d076d065b00360bb201af0ba1046a074301b60c3308b50a45068305040c5a017f057d0322013101ea04680bbf01b60b2f08ce08ad05490c1801b10aec04230809003902e107840219068207b5029c032a0b8c01d40cfd09a7054707f10aca0c03081e0cf502800843050506c100aa0ac707c7054e03ba05bf0a29065603d60c2107b005a1080e097201740b9409bd0ce20b9f00b8077b01020a590c0509ca09960a48011e0430020708eb067a04b70c0b0bde01a9070a068d0c180a0b07a60bcc0c3d023b092005e80aa004db01ec057a061807af04f8020b09fe05050a5f00d90c8f0af5064e087d067b09b302a30567
5.04740aed04500b5a062b022b069907ac030b0c530696068d07880c7d041f06dd0a5c0b650c0e0534082c054a05800bf90abf016801e605e906a3067f098500a6019e0bf6062c04080ba70b190123004106dc01e4069b01db04d9056f0ab5055306300ca0014800e80204074f0ce707f2009d09220816066a09350751068408be063a01b9053a033d08320148019e0b3e0b26039007f808e80177090805ec019c08ea08cb06b3026d0332029506f3014802780799099d01f602150494047c07b308200a25046303e708bf0897082c035503b4051b06110b890c3900430afc08aa07aa075f0674058c0a8a028f012e089a077902440c020b870a38022801c2098406c101e70651031e003d037705760ab6053c073b0a9109a004750a550221058507a806f1021d0c67091602300845020f01d207a605b3019d0a980195062c0ac10bdb06fa01a3077d0054088400540c5709710c48022a045202590635013501080bcf04020b3f057d067c09c5003002170b0b0499062607af00d8075d0aed0a3503bb0a840c04044c05520ad4080f09c40b1b08df009c00990afc04160b82036f0b4309c90566004b007408d508e509990a530af306910cd30499029b0a4f05370c700677032103ec0c8304e0012e053505a50567098705c70ae2064a09da05cf00e9054a054707510c4a00d7019c04750ba60c8706f30c89076908cc09d50693
6.061303b608940614076e01eb0cd90aca08a20544087902e803f5074c02f20bed09d909e0031104f807ce092606550a5405be01ef015a0a95080304e2027207410c9905c20c79003d0c710c0c071d05c70312031f00d004a0016c043d0001048f03f506b50cff0871066208b40a5d075a0b4c09700865065102cc07170a790972019c06b80a860a280b92067306c90b050a3e0b77014903e0005e01bc0a7a0b0f021b077b024d08290ca50a7d015402c1087e068500810b6e024c05a1011d03a2035c0b7b0c62062d0b9d069102630cd00b1f08cc05b30c9c008603280aa203300b1105aa000d0cb40c870cc602bb020707670cd007140ad602200aa90ae604510958060104de0b620164047d092e06d60050049b080903460c21056301ca056f0b3807b600bf051401ca094909f60bf40cf106be039605180a700a0f04b50a410a0e08a0084c08db07cf01d1029106d7055a0048043c0c78009500f9052c082f0bca030a050e0200013d0993020c09df0264036a06cb02140a9d03b30b9a09ba0310080e0cb90a2c075407c7045606a90ac004f509d0046a0ba30bb50aef072e07a0071e06f009240664017d0c0e0b440ce206f50b960ae80238023e03050aeb0c6b09dd008d05ac0459035403b30765045208f002eb04d106390aed0a5405f500c9021a04ed0cb601e704980a720c6b07c109ef01f301c409490011007f0a6b
7.04ea01ef047504e1023f056e080f0bff0b7e0b4b0c0108460179064203ea01e009b10033039c01d109fa03ef01660184082907bc099c099802fa02c8016c08ae0b110a6d0711007a067c07690173084d0a54028d030f045804cb0038044b0bf006bb006104b90a2d0ad708f808a40ce903b7019d0c530a5605cf01b407d80c1c047a0c4d02bb095d016e061706af07a208c104430bdf08120c39021401aa022a029907bf07b700ba09a90a0e055a05f20aa4048501c901810add01470be90c88092707d609d203030a7a021e089f0cc5061d05c8027707c1089707540af106e10c8e036c04d5094504720075090f03c208ea0b3f00e60b01061e02ec0a3f08f9051e01c6063d0972097801f7095404f7059c088e03a200d3081105ef03850b5a0960090b06f903e8042002bb07470bcd0456016b01910bdc0be800a901330598085f014908b60bfc003307b8045002a501800cf703f80665030805d90298018c0b9f02fc094707d4031d01e90476042801f008840b7f0ad805fc02e405ce0729024c056104cd044106090cde01380c5f07b8047c07b50b4c03400bbf02b901c1081908420c43098707bc01e102e5042805c80150040805ad05580b3f0398027e05e90c7b01d40307041a0b9501c60be9014300ff0002028b0470013508520a76043d047901050a6d009309810a95044c069c046c04a3002a07ff06430b5103ea
8.03dd01930a1605e90800076903fb07c7056a079c085d035e031c06890011054206030c9f019408400791027e00c10c4e054008840b6c007809f20c8700fb034b03480c010cf703410672001f06520cbc021d0786070e052c047a0c990b4c056e017b028e004e0a390972007d0b2d0660066c0324009c0a96084a0c480a370ce000160644077a029e066800a60a02012a0a6a05630a6e0281049f01b2047f068e08780529043d07c604d6027d0b3e0b9d0611043404a1046209ac050705f6096c0b7f00e802570798055e03770989076f08010b0204e304cd081c017c070503150bc202c201fc048403230cd60b8802a0005d074003a801de081407d802990cce0a2806b40b1f0743042e005302b80ab2048502220a590bd903e70230007f0ad804bc0a020c1b01f70cf6045e021f00910c0c048a019d09df0c3703c6096305fe010c0bef0790017f072a0588065f03f3003a0a2701c8045403d008f20bdc042d02ee0c4e09ec034a02710ab40b2103f00434093f090d031f055c029507d50c39019e0a19069506e00533038a040d090a08780b15004504490350017700fb01d3032c07bf09010a4603bd040800ff0cc2084f04da06e4039401800c75082308890411008e099f08880aa60ae4057707bf0c240403021306ca074c096908d1093409db003809da02c70845069404ef06ad096303fe0a7500b907e60c5004660caf
9.003000ac09cb0bb4030501e8042a061c065f05d200710a2d07630042062c03620b77003007d90447067800b509b403d100a1043c0a23050a09ec0b1a06790a1809a702300cce0596051701dc05b108e20844096f06ac0862005209be006700540a7f0103009705b30a81081c05e6092e09050491036302db02c40a620050047601ed04fb02fe002d0cbf01240a020a0a0ca7040101e501760b7b0047089f011a0cd60a3808ea0c9d0666052b0306091307cf015107ae0419079407a20b7605ad03bb09b90b06078e056602c00c440996072c012703a3082600f0001f00ad048c01ea04fe0af50541084307e30a2c0b36036a0cb509310d000b1406cf00550a800ae908ff0a2704b209a1006f049906c4076304a20a140b5803b207be04570842089203410050045f053207f70377005b01b0006b0acc08150233078a0be509a20af70b66065a070e0cd00c62064b0569044a0594056d08b705fa052900b8070d072f09ea0645090200b60069006d09f7043003e7059f06d502f9019107f207df04890063074b0c3707270c5c0a18023802b406f80ce30541083e0b1008cd01a10bfc024609f10a75078e03e40ab008e9082d0a5e0a1609200c4404fd047b08910092020f09360af10add0c21004409ff09f802b400120755047906fe050205e706cf01aa0c4504da03f804470b950005032a03c703ee052307de05080086007f
*/

/*
Public Matrix Poly 3x3 (coeff 0 -> coeff 256), 16 bits per coef
public matrix poly 0: 06db059e0a360c1f05db08780c010a9200df0cb902330ca9003400e00a5f0adb054c076f06620249098803d10731022308ca059307130983009f02d5089109af0b9b0b4706d2055c09480b8a075b022c0487043f0a2500bd0378008700540c2d050e0b9500e9024a0687093b052903a90a7e00da0636014a0bb206840036086a06600cb902780840064b06c8079a01f00595069c067800b20bd30c850bdc07f40c3d02e709df053c072d0794071f04af042f085d019a089b0a9e0443024001ce079d047901aa0c340aca00f904400a8b01b908da06ff0cb50c22072603f303a50ba201ea054604d605fd01300b7c0cb10714037e09d80a1a08b401f504450cf400dd058e0912023e0c48029e02620acd0c2d0b7a06e40aa30432080203c707ca083704d50ab60b6f0888003203b000150a5d08af06c70496026b0229014202a00a8a04c201050ac1077106640c2909df015809370892080709ed09c0035f06490c4e09b7006207e303a7087309ae0ca608c704d904480c2b064c0b0e098a044b0a7d014c0aa6003204250b71069305f3032e0c15068201d0080200c10ca7059901a90a7401780059011206d900e30408090500ce081909f102f206a80094067a02ac01a00b16045302d9045703000250063608d6075903130a7903d901f8030b08d305160a3b0183066400230732043709b20813051706d6024708c40ce501ae
public matrix poly 1: 07f20947066405770c060c1002090c0407bd0c0706900ab00bbc00df071001fb04b007fd0ce9086d068204b3058400400093058f0ca900c901e606070be2069804b80b6809500cae0aa1041e037c038105820ac3084c0c26040f0b720ab306ed0d000aed0bb50a7a01980bf40c560a7f0cea0bd90c8409590b8b091a02650c2f08ee06150c5800230cd008a10a71086203df01a20a78047000320b680c560ac409e70ccc0544081e095a09300100081505fc017304fa08f904b004ad09d5053401dd061308230409051e0121037e08cf011200f5054a066c048d070c07df031a007701e30431024c08aa04bb0b93078a01e9090e05c50cbc015608ee03660b6100da057200f30c1a07030bac0cb1019e01ea0292052804b5028f0b8906bf00b007f602270a750954014501d503b403db0369048a069106b902ac08230a800909061305680b3402d60bb706420a8d05a20a9c08d903e80c370bbb033706c10a8a0a980b7e0486080003c800300c9f026d057004b7067c08460a0b0117061f00ce051603af05d60a1b084a07c4077a03680ca407fa0c4206a0086300ac0bd90c4b015808ee03f30b2e011d003e0a14004209e90b4d0624050d057e039d03e400aa04a205b102710cab0be6050f0d0005e20188064e0761023d057f0a5901fa011709ca0108017c052b08b90aae0bc8021903da0c61002f0cd40276037609f406dc
public matrix poly 2: 08a70cd402fd05b606570562017706a30406045206ea098a01ab0a9d0ad9034f0560033506ed094a09c5088b074f05e503ee0c0a0076016f0a2e04b400c00100013a039b0c640b8e00b8084d0c92023a066902f4051303b30b6d050b014c068605d30723014c00960c910431026c02db094e0508056e050c07a60a590a0f04020a3f059f01f607530161029a009602e90c3f01f6072602bf0aad01f5060403300cfc03ff01c301f001f309f004be0128044f098908b70727000a076601bc0b3f00e808c10a9f0c6504ed03b904120a7d07ba0aea004e0aad0ab40c8807f90c9707ce064600270745005005670ba3003b06f403e00a5f05b10c11055b06ee06c1035808b303c20ae90c560be7095a081e0b800a80049f015c0ca200520509026e0752071e08c001730460033007d20b15088a0a5a0b590bcb06200480044700e609430c5c0bef0be608c9027b063a0b55081603c8036b06da0704064407e103b001320b1e05fa07f203f000e407bc00cf03020511025903ec036105f100c902c4047505fe0c1a00200530036d0ade01aa09e60baa072d090700a906af08eb075407bb040e0632046c05ed0cd3081705d000c00c3404ea03ce0b37009b0c5804b3076f0876099c05cf0aac081007fe0b270b700a6007000182098500170c390545083b07da0c1b01d10b0c050c0cdb022a0ab60772043604080497088305df04d4
public matrix poly 3: 056702a309b3067b087d064e0af50c8f00d90a5f050509fe020b04f807af0618057a01ec04db0aa005e80920023b0c3d0bcc07a60a0b0c18068d070a01a90bde0c0b04b7067a08eb02070430011e0a48099609ca0c050a590102077b00b80b9f0ce209bd0b9401740972080e05a107b00c2103d606560a2905bf03ba054e07c70ac700aa06c10505084302800cf5081e0c030aca07f1054709a70cfd01d40b8c032a029c07b506820219078402e10039080904230aec01b10c18054908ad08ce0b2f01b60bbf046801ea01310322057d017f0c5a050406830a4508b50c3301b60743046a0ba101af0bb20036065b076d013d02cc04ce001e08200c76007100fd00390c55084505bb0b6e0a540733089a072805410312049403cb0a1106bc03d1047507f700060aa601ef00d605710cfc00020c8e04bb002307b20848072b0c66089c040a0c0803e0001c041b028d04ee0592039605f10aba0027032007fe004c047708540810051a02a60c630ac906a90a0e039d049408dc01a706430b31019903e508f00aa20860041002c301fb087e01140c000cac09cb08540c96080d04ec01fd099906a80774018302840a59021207b4097405e504970b8c09af0a2605ce09600b540b4c08ab07c50844000e0646015b04a102e900ef0684096a09f202540ade0bbb097f05ea0c070a4e0b4b0beb0a830968007b05f40529068e0c9901a4
public matrix poly 4: 069309d508cc07690c8906f30c870ba60475019c00d70c4a07510547054a00e905cf09da064a0ae205c70987056705a50535012e04e00c8303ec032106770c7005370a4f029b04990cd306910af30a53099908e508d50074004b056609c90b43036f0b8204160afc0099009c08df0b1b09c4080f0ad40552044c0c040a8403bb0a350aed075d00d807af062604990b0b0217003009c5067c057d0b3f04020bcf01080135063502590452022a0c4809710c57005408840054077d01a306fa0bdb0ac1062c01950a98019d05b307a601d2020f0845023009160c67021d06f107a8058502210a55047509a00a91073b053c0ab605760377003d031e065101e706c1098401c202280a380b870c0202440779089a012e028f0a8a058c0674075f07aa08aa0afc00430c390b890611051b03b40355082c089708bf03e704630a25082007b3047c0494021501f6099d07990278014806f302950332026d06b308cb08ea019c05ec0908017708e807f803900b260b3e019e01480832033d053a01b9063a08be068407510935066a08160922009d07f20ce7074f020400e801480ca0063005530ab5056f04d901db069b01e406dc004101230b190ba70408062c0bf6019e00a60985067f06a305e901e601680abf0bf90580054a082c05340c0e0b650a5c06dd041f0c7d0788068d06960c53030b07ac0699022b062b0b5a04500aed0474
public matrix poly 5: 0a6b007f0011094901c401f309ef07c10c6b0a72049801e70cb604ed021a00c905f50a540aed063904d102eb08f00452076503b30354045905ac008d09dd0c6b0aeb0305023e02380ae80b9606f50ce20b440c0e017d0664092406f0071e07a0072e0aef0bb50ba3046a09d004f50ac006a9045607c707540a2c0cb9080e031009ba0b9a03b30a9d021406cb036a026409df020c0993013d0200050e030a0bca082f052c00f900950c78043c0048055a06d7029101d107cf08db084c08a00a0e0a4104b50a0f0a700518039606be0cf10bf409f6094901ca051400bf07b60b38056f01ca05630c2103460809049b005006d6092e047d01640b6204de0601095804510ae60aa902200ad607140cd00767020702bb0cc60c870cb4000d05aa0b1103300aa2032800860c9c05b308cc0b1f0cd0026306910b9d062d0c620b7b035c03a2011d05a1024c0b6e00810685087e02c101540a7d0ca50829024d077b021b0b0f0a7a01bc005e03e001490b770a3e0b0506c906730b920a280a8606b8019c09720a79071702cc0651086509700b4c075a0a5d08b4066208710cff06b503f5048f0001043d016c04a000d0031f031205c7071d0c0c0c71003d0c7905c20c990741027204e208030a95015a01ef05be0a540655092607ce04f8031109e009d90bed02f2074c03f502e80879054408a20aca0cd901eb076e0614089403b60613
public matrix poly 6: 03ea0b51064307ff002a04a3046c069c044c0a95098100930a6d01050479043d0a76085201350470028b000200ff01430be901c60b95041a030701d40c7b05e9027e03980b3f055805ad0408015005c8042802e501e107bc09870c430842081901c102b90bbf03400b4c07b5047c07b80c5f01380cde0609044104cd0561024c072905ce02e405fc0ad80b7f088401f00428047601e9031d07d4094702fc0b9f018c029805d90308066503f80cf7018002a5045007b800330bfc08b60149085f0598013300a90be80bdc0191016b04560bcd074702bb042003e806f9090b09600b5a038505ef081100d303a2088e059c04f7095401f709780972063d01c6051e08f90a3f02ec061e0b0100e60b3f08ea03c2090f00750472094504d5036c0c8e06e10af10754089707c1027705c8061d0cc5089f021e0a7a030309d207d609270c880be901470add018101c904850aa405f2055a0a0e09a900ba07b707bf0299022a01aa02140c3908120bdf044308c107a206af0617016e095d02bb0c4d047a0c1c07d801b405cf0a560c53019d03b70ce908a408f80ad70a2d04b9006106bb0bf0044b003804cb0458030f028d0a54084d01730769067c007a07110a6d0b1108ae016c02c802fa0998099c07bc08290184016603ef09fa01d1039c003309b101e003ea0642017908460c010b4b0b7e0bff080f056e023f04e1047501ef04ea
public matrix poly 7: 0caf04660c5007e600b90a7503fe096306ad04ef0694084502c709da003809db093408d10969074c06ca021304030c2407bf05770ae40aa60888099f008e0411088908230c750180039406e404da084f0cc200ff040803bd0a46090107bf032c01d300fb01770350044900450b150878090a040d038a053306e006950a19019e0c3907d50295055c031f090d093f043403f00b210ab40271034a09ec0c4e02ee042d0bdc08f203d0045401c80a27003a03f3065f0588072a017f07900bef010c05fe096303c60c3709df019d048a0c0c0091021f045e0cf601f70c1b0a0204bc0ad8007f023003e70bd90a59022204850ab202b80053042e07430b1f06b40a280cce029907d8081401de03a80740005d02a00b880cd60323048401fc02c20bc203150705017c081c04cd04e30b020801076f09890377055e0798025700e80b7f096c05f6050709ac046204a1043406110b9d0b3e027d04d607c6043d05290878068e047f01b2049f02810a6e05630a6a012a0a0200a60668029e077a064400160ce00a370c48084a0a96009c0324066c06600b2d007d09720a39004e028e017b056e0b4c0c99047a052c070e0786021d0cbc0652001f067203410cf70c010348034b00fb0c8709f200780b6c088405400c4e00c1027e0791084001940c9f0603054200110689031c035e085d079c056a07c703fb0769080005e90a16019303dd
public matrix poly 8: 007f0086050807de052303ee03c7032a00050b95044703f804da0c4501aa06cf05e7050206fe04790755001202b409f809ff00440c210add0af10936020f00920891047b04fd0c4409200a160a5e082d08e90ab003e4078e0a7509f102460bfc01a108cd0b10083e05410ce306f802b402380a180c5c07270c37074b0063048907df07f2019102f906d5059f03e7043009f7006d006900b60902064509ea072f070d00b8052905fa08b7056d0594044a0569064b0c620cd0070e065a0b660af709a20be5078a023308150acc006b01b0005b037707f70532045f0050034108920842045707be03b20b580a1404a2076306c40499006f09a104b20a2708ff0ae90a80005506cf0b140d0009310cb5036a0b360a2c07e3084305410af504fe01ea048c00ad001f00f0082603a30127072c09960c4402c00566078e0b0609b903bb05ad0b7607a20794041907ae015107cf09130306052b06660c9d08ea0a380cd6011a089f00470b7b017601e504010ca70a0a0a0201240cbf002d02fe04fb01ed047600500a6202c402db036304910905092e05e6081c0a8105b3009701030a7f0054006709be0052086206ac096f084408e205b101dc051705960cce023009a70a1806790b1a09ec050a0a23043c00a103d109b400b50678044707d900300b770362062c004207630a2d007105d2065f061c042a01e803050bb409cb00ac0030
*/

// Comparing SHAKE output with C (4032 bits)
// poly 1:9d9747aa41c3ca9a0f40b4a8c79e1bdaf86fb52cc226373fa523bab2af1e46e5fd046f4dfd05137d5dde7c1bcb584e717e93d03e8f9d1a4a8bf581f7455d44f4dc0d8e25913e82c417ef29bf2d26cddac2c9adb74efeeee4e6d3f13faaa12e430258e5c7a37c37584db6fab6008f8832003b15d0a5af18dcc766496b922242012a8a2a4c0511ac71476629fc9d5871939278803bdf9ec049e75f83da4956fc4e7c9b62307e6ffdf1a73387ae69ca267e8cd9844473bfc24ce6b08ab9447dca14a62a032514b71a3d69f3e532152c68d02180c170ca99951a748a17592011d946dbe3e0d14d8e4005e90c19189ff2826a94a067ac021ac76db1699ee2b6ddda083f45e29e2d537e4500032536668d5917fb1c4fe8a73f31799a3df8b130d368513b3a18a24f6623207337249b137851d67624c458ce6cef1a63257e3d92cb61cce10f9e979049a6d9b3194fcaa2f5743b976a9de7b4dcf61568e639cf61df867ba391d6f27bca44f5adac07e09e088cda63f8a5214450ce313e350c10a65d34975041a73f78c8968c6e75a0895adc506359095ccdb936cbbf2426fb53fdc53414cddeb8d6a95de8a9debd8634ebeb861ca0d3551feef5f4b39154acb90c697ec1d25101950fac0623a53fef8647ce485b07a082e9c2d7dd598b053984b21916ee66a153528fb631255541f9b4e5ae8fe837a706c2ced50679