../params.vh