`timescale 1ns / 1ps
`define DELAY 3
// for noise, gen e1,e2,r in kyber768
// e1, r = output poly 3 times (1024 bits each)
// e2 = output poly 1 time
// for public matrix, gen A transpose (9 polys)
// run once, collect 7 polys?
module hash_top_tb;
  reg clk;
  reg enable;
  reg rst;
  reg [255:0] coins;
  reg [255:0] seed;
  reg [3:0] domain;
  reg [13:0] output_len;
  //// output
  wire [4095:0] noise_poly_out;
  wire [4095:0] public_matrix_poly_out;
  wire noise_done;
  wire public_matrix_done;
  integer i;

  hash_top hash_top_uut (
        .clk(clk),
        .enable(enable),
        .rst(rst),
        .coins(coins),
        .seed(seed),
        .noise_done(noise_done),
        .public_matrix_done(public_matrix_done),
        .noise_poly_out(noise_poly_out),
        .public_matrix_poly_out(public_matrix_poly_out)
  );
  // reverse bytes for printing (this time, per 4 bytes)
task print_decimal_pm(input [4095:0] S);
    integer b;
    localparam integer NUM_BYTES = 256;
    //reg [4095:0] reverse_coef;
    logic [15:0] coeff;
    begin
        // reverse bytes (for visualization)
        for (b = 0; b < NUM_BYTES; b = b + 1) begin
            coeff = S[16*b +: 16];
            // print as deci
            $write("%0d ", coeff);
        end
    end
endtask

  initial begin
    $dumpfile("dump.vcd");
    $dumpvars(0, hash_top_tb);
    clk = 0;
    forever #(`DELAY / 2) clk = ~clk;
  end

 initial begin
    // -- INPUT -- //
    rst = 1;
    coins  = 256'hf8f11229044dfea54ddc214aaa439e7ea06b9b4ede8a3e3f6dfef500c9665598;
    seed = 256'hf8f11229044dfea54ddc214aaa439e7ea06b9b4ede8a3e3f6dfef500c9665598;
    enable = 0;

    // Release reset to start loading state_reg, done, etc
    #(`DELAY) rst = 0;
    #(`DELAY) enable = 1;

    wait (noise_done == 1'b1);
    wait (public_matrix_done == 1'b1);

    #(`DELAY * 5);

    $display("\n\nnoise output from SHAKE : %h\n",hash_top_uut.noise_stream[1023:0]);
    //print_state_bytes(hash_top_uut.noise_stream[1023:0]);
    $display("\n\ndone : %b\n noise string (4096 bits) = %h\n", noise_done, noise_poly_out);

    $display("CBD coeffs (0..255):");
    for (i = 0; i < 256; i=i+1) begin
        $write("%0d ", $signed(noise_poly_out[i*16 +: 16]));
        //if(i%16==0 && i!=0) $display();
    end

    $display("\n\npublic matrix output from SHAKE : %h\n",hash_top_uut.public_matrix_stream[5375:0]);
    //print_state_bytes(hash_top_uut.public_matrix_stream[5375:0]);
    $display("\n\ndone : %b\n public matrix string (4096 bits) = %h\n", public_matrix_done, public_matrix_poly_out);
    print_decimal_pm(public_matrix_poly_out);
    wait (public_matrix_done == 1'b1);
        @(posedge clk);  // +1 clock
    $finish;
 end
endmodule

// CHECKING PUBLIC MATRIX OUTPUT
// Public Matrix from SHAKE : b17a22ce5d458ba33d6931d893324e04123b1590846653d49d019a59da9ddd1aad293fc43863b0f63c093b2e9325249a0e45cf390f8ea91fdf9450a90c34babde106958e80184c9dfcf78da5f66fd7f65feef73aced58d4d995606c2ab56d11141ec5e47c6c8baaa5fcc346f9ea76c58389af2cf4df93f38c70f542cbae644577d22fd10d46f4f5c70d72c99775bc9ed7e0c417b6af0e9e545603f42df15d09481539cfef0bdb84b3899339793c2759f4c6d3b73f07f5a2ef7927f39a6ca2b45102a5b2794449c99b04617b2bee4777e043007a9e07eb858f4a49fdb5380e1de3b739c795715f4fc11223f37896d5fce01f63ce25780c462a6f9379a8d112d026133e5b6b6df3795cc374c51785f435d2bcf64e4f6be21e38f7d8c1c447b2e73b9ca12d58a71efbc7d4cae4cb99541d8f5662dc2ad1b4083c449461b60e7ca6bd395bc878cd37eff6ebca7ec10ee6ffbe1f719eec9ebbfd31e60b174c4e4a2940d14ce9343b3c10d9ddd42d92d04c19c1ae1901cb4095fa4e00ee14949ad2f513257e1bc6295e8a0eda314c3ac3b67a0d62a4397efedd96eed0ecba9cc195276800fa0bd99a52dcdbe8d959276e5ace0fb215f3a7b01d781ef77287786653a6e7a15c187709b16854e142910976b0987ac13fd54981c47af0635eb286caeadd9c25c425088160c7965659c1e659c9a5942b330dd5f045ddf6689eac9ea06a1bd59b27768331e8b8d74f8b5c661789989160286a71e740bcd0718d5e8b84a05bdb9aa0964512c452e2feec81ad94069ce5430a05d5b806d311a9a913492a419012859b1884f94698c62a85ac0d7cf91e370d3a14a0d75d1ee3177b29cdf4aac5463b73d722603fcd1c946b71f4d60b1d0619be63b2c10464e8eed2db46d0fa6ba16beaa63a2f5f9ff6ccbe3e70953c633e81da07d3389ef6becfcfdba740b56bc
// After Sampling Rejection : 07100291044e0851069b070807c101570a6e03a605860772087701d700170b3a05f201fb0ce50769029508db02da05990bda000f08070652019c0ca90cb006ed09ed074302ad06a006730bac0c3104a300e8095602bc07320512049409e100ee00a405f009b401c900e101a90cc10042042d00dc01b3043903ce01400a2e04c4074b016001ed03bf09ee019f07e1010e0ca70bc607ed038c087b0c950bca001b046409c40834001b0adc022d066f05d8041905b904ca07db0cef07180ad5012c0ab9073204410c8c07d8021b04cf02b505f7085104c307cc095307df0b6b06e50336010202d1018d09a307f90a6602c4080507e203cf06010ce50893073f022101fc055707990c7303bd080503db09fa04f4058b087e09070300047e077e04be0b2107460b09099c0449042705b20a1004520bca0a63097f092f072e05a707330b6d04c90c2903970339093804bb08bd0538019405df0423045e05e90a7b04100c7e095b0779092c005c04f6010f07d507440a2c0540038304dc09a3085806ca079e06f304cc05fa0aba0c8c064705ee0c41011d01560abc02060569094d08dd05ce03af07ee05ff06d706ff06a508df07fc09d40c180808006e01bd0ba3040c0a95009408e00cf4050e09a20425093200930cf60b0603380c430ad10add09dd0a5909a0019d03660849001503b1020404e30293016903da038b045502270ab1
// Reverse coeffs to compare with C : 0ab102270455038b03da0169029304e3020403b1001508490366019d09a00a5909dd0add0ad10c4303380b060cf600930932042509a2050e0cf408e000940a95040c0ba301bd006e08080c1809d407fc08df06a506ff06d705ff07ee03af05ce08dd094d056902060abc0156011d0c4105ee06470c8c0aba05fa04cc06f3079e06ca085809a304dc038305400a2c074407d5010f04f6005c092c0779095b0c7e04100a7b05e9045e042305df0194053808bd04bb0938033903970c2904c90b6d073305a7072e092f097f0a630bca04520a1005b204270449099c0b0907460b2104be077e047e03000907087e058b04f409fa03db080503bd0c730799055701fc0221073f08930ce5060103cf07e2080502c40a6607f909a3018d02d10102033606e50b6b07df095307cc04c3085105f702b504cf021b07d80c8c044107320ab9012c0ad507180cef07db04ca05b9041905d8066f022d0adc001b083409c40464001b0bca0c95087b038c07ed0bc60ca7010e07e1019f09ee03bf01ed0160074b04c40a2e014003ce043901b300dc042d00420cc101a900e101c909b405f000a400ee09e104940512073202bc095600e804a30c310bac067306a002ad074309ed06ed0cb00ca9019c06520807000f0bda059902da08db029507690ce501fb05f20b3a001701d708770772058603a60a6e015707c10708069b0851044e02910710
// Coef from LSB to MSB order : 2737 551 1109 907 986 361 659 1251 516 945 21 2121 870 413 2464 2649 2525 2781 2769 3139 824 2822 3318 147 2354 1061 2466 1294 3316 2272 148 2709 1036 2979 445 110 2056 3096 2516 2044 2271 1701 1791 1751 1535 2030 943 1486 2269 2381 1385 518 2748 342 285 3137 1518 1607 3212 2746 1530 1228 1779 1950 1738 2136 2467 1244 899 1344 2604 1860 2005 271 1270 92 2348 1913 2395 3198 1040 2683 1513 1118 1059 1503 404 1336 2237 1211 2360 825 919 3113 1225 2925 1843 1447 1838 2351 2431 2659 3018 1106 2576 1458 1063 1097 2460 2825 1862 2849 1214 1918 1150 768 2311 2174 1419 1268 2554 987 2053 957 3187 1945 1367 508 545 1855 2195 3301 1537 975 2018 2053 708 2662 2041 2467 397 721 258 822 1765 2923 2015 2387 1996 1219 2129 1527 693 1231 539 2008 3212 1089 1842 2745 300 2773 1816 3311 2011 1226 1465 1049 1496 1647 557 2780 27 2100 2500 1124 27 3018 3221 2171 908 2029 3014 3239 270 2017 415 2542 959 493 352 1867 1220 2606 320 974 1081 435 220 1069 66 3265 425 225 457 2484 1520 164 238 2529 1172 1298 1842 700 2390 232 1187 3121 2988 1651 1696 685 1859 2541 1773 3248 3241 412 1618 2055 15 3034 1433 730 2267 661 1897 3301 507 1522 2874 23 471 2167 1906 1414 934 2670 343 1985 1800 1691 2129 1102 657 1808
// From C official : 2737 551 1109 907 986 361 659 1251 516 945 21 2121 870 413 2464 2649 2525 2781 2769 3139 824 2822 3318 147 2354 1061 2466 1294 3316 2272 148 2709 1036 2979 445 110 2056 3096 2516 2044 2271 1701 1791 1751 1535 2030 943 1486 2269 2381 1385 518 2748 342 285 3137 1518 1607 3212 2746 1530 1228 1779 1950 1738 2136 2467 1244 899 1344 2604 1860 2005 271 1270 92 2348 1913 2395 3198 1040 2683 1513 1118 1059 1503 404 1336 2237 1211 2360 825 919 3113 1225 2925 1843 1447 1838 2351 2431 2659 3018 1106 2576 1458 1063 1097 2460 2825 1862 2849 1214 1918 1150 768 2311 2174 1419 1268 2554 987 2053 957 3187 1945 1367 508 545 1855 2195 3301 1537 975 2018 2053 708 2662 2041 2467 397 721 258 822 1765 2923 2015 2387 1996 1219 2129 1527 693 1231 539 2008 3212 1089 1842 2745 300 2773 1816 3311 2011 1226 1465 1049 1496 1647 557 2780 27 2100 2500 1124 27 3018 3221 2171 908 2029 3014 3239 270 2017 415 2542 959 493 352 1867 1220 2606 320 974 1081 435 220 1069 66 3265 425 225 457 2484 1520 164 238 2529 1172 1298 1842 700 2390 232 1187 3121 2988 1651 1696 685 1859 2541 1773 3248 3241 412 1618 2055 15 3034 1433 730 2267 661 1897 3301 507 1522 2874 23 471 2167 1906 1414 934 2670 343 1985 1800 1691 2129 1102 657 1808
// Reverse Sampling Verfied : 16/1/26

// CHECKING NOISE OUTPUT
// Noise from SHAKE : 99abf40515a7387aa7a41f83840467aaba58818583cae85ec7710efbeb5dce0a5e91f3fa854b8570aaa4393e663ef90458d0d9823e682c1062947b54c496ef8a9bb38198777295bb264c790628226b8a3a3ce2172d0d0c5534d8dc67d0c1155c4a98b3559c84fa82d90e4cfc474b2fda6b38ca4f0ef964bd4efd4b5cd5be6696
// After cbd :  00000000000000000001ffffffff00000000fffeffff00010000ffffffffffff0001ffff0000ffff000000000000ffffffff0000fffe00000002ffff00000001ffff000000010000ffff0001ffff00010000fffefffffffe0000ffffffff0000ffff000100000000ffffffff0000fffe00000000000100020000ffffffff00000000fffe00010000fffe0001ffff000000000001fffffffeffffffff0002ffff000000000000fffe0000ffff0001ffff00010001ffff00010002fffe00020000ffff000000000001000100010001ffff0000000000010000fffffffe00010000000100010000000000010001000100010000ffffffff00010001000200000001ffff0000ffff000000000000fffeffff0000ffff000100010000ffff00000001000100000001fffe0000ffff0002ffffffff0001ffff0000ffff00000000ffff0000ffff000000000002ffff000000000002ffff000200000000ffff0000000000010000ffff0000ffff0001ffff00000000000000000002000000010000ffff00000000fffeffff0000ffffffff0001000000010000ffff00010001fffe00010000fffffffffffffffe0000ffff0002ffff0000ffff00010000ffff0001000000000000000000010000ffffffffffffffff0002000100000000ffff00000001000100000002ffff0000000100010000000000000000ffff0000000100000000
// Coef from LSB to MSB order : 0 0 1 0 -1 0 0 0 0 1 1 0 -1 2 0 1 1 0 -1 0 0 1 2 -1 -1 -1 -1 0 1 0 0 0 0 1 -1 0 1 -1 0 -1 2 -1 0 -2 -1 -1 -1 0 1 -2 1 1 -1 0 1 0 1 -1 -1 0 -1 -2 0 0 -1 0 1 0 2 0 0 0 0 -1 1 -1 0 -1 0 1 0 0 -1 0 0 2 -1 2 0 0 -1 2 0 0 -1 0 -1 0 0 -1 0 -1 1 -1 -1 2 -1 0 -2 1 0 1 1 0 -1 0 1 1 -1 0 -1 -2 0 0 0 -1 0 -1 1 0 2 1 1 -1 -1 0 1 1 1 1 0 0 1 1 0 1 -2 -1 0 1 0 0 -1 1 1 1 1 0 0 -1 0 2 -2 2 1 -1 1 1 -1 1 -1 0 -2 0 0 0 -1 2 -1 -1 -2 -1 1 0 0 -1 1 -2 0 1 -2 0 0 -1 -1 0 2 1 0 0 -2 0 -1 -1 0 0 1 -1 0 -1 -1 0 -2 -1 -2 0 1 -1 1 -1 0 1 0 -1 1 0 -1 2 0 -2 0 -1 -1 0 0 0 -1 0 -1 1 -1 -1 -1 0 1 -1 -2 0 0 -1 -1 1 0 0 0 0 
// From C official : 0 0 1 0 -1 0 0 0 0 1 1 0 -1 2 0 1 1 0 -1 0 0 1 2 -1 -1 -1 -1 0 1 0 0 0 0 1 -1 0 1 -1 0 -1 2 -1 0 -2 -1 -1 -1 0 1 -2 1 1 -1 0 1 0 1 -1 -1 0 -1 -2 0 0 -1 0 1 0 2 0 0 0 0 -1 1 -1 0 -1 0 1 0 0 -1 0 0 2 -1 2 0 0 -1 2 0 0 -1 0 -1 0 0 -1 0 -1 1 -1 -1 2 -1 0 -2 1 0 1 1 0 -1 0 1 1 -1 0 -1 -2 0 0 0 -1 0 -1 1 0 2 1 1 -1 -1 0 1 1 1 1 0 0 1 1 0 1 -2 -1 0 1 0 0 -1 1 1 1 1 0 0 -1 0 2 -2 2 1 -1 1 1 -1 1 -1 0 -2 0 0 0 -1 2 -1 -1 -2 -1 1 0 0 -1 1 -2 0 1 -2 0 0 -1 -1 0 2 1 0 0 -2 0 -1 -1 0 0 1 -1 0 -1 -1 0 -2 -1 -2 0 1 -1 1 -1 0 1 0 -1 1 0 -1 2 0 -2 0 -1 -1 0 0 0 -1 0 -1 1 -1 -1 -1 0 1 -1 -2 0 0 -1 -1 1 0 0 0 0
// CBD verified : 16/1/26