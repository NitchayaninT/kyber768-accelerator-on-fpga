`include "params.vh"
module polyvec_pointwise_acc_montgomery (
  input [15:0] a [256][3],
  input [15:0] b [256][3],
  output [15:0] r [256]
  );

  reg [5:0] i;
  
endmodule
