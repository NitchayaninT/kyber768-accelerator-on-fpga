package params_pkg;
  parameter int KYBER_K = 3;
  parameter int KYBER_N = 256;
  parameter int KYBER_Q = 3329;
  // ... other parameters
endpackage
