module rho_tb;


