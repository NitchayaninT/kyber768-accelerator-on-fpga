module poly_basemul_montgomery(
  input [15:0] a [255],
  input [15:0] b [255],
  input clk,enable,
  output [15:0] r [255]
);

  reg [5:0] i;

  always begin
  end
endmodule
