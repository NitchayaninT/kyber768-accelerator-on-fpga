`timescale 1ns / 1ps
`include "params.vh"

// each coefficient in polynomial ring use on cla_adder
// 4rounds of addition is made and then copy value from buffer to output
